LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY projetoelevador IS
PORT ( SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		LEDR : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		display: out std_LOGIC_VECTOR(6 DOWNTO 0));
END projetoelevador;
ARCHITECTURE Behavior OF projetoelevador IS
BEGIN
LEDR <= SW;

Case SW is
	when SW(1):='1' <= display <= "0000001";



END Behavior;